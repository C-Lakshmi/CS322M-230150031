// NOT gate
module MyNot(input A, output Z);
  assign Z = ~A;
endmodule
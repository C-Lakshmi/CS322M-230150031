// AND gate
module MyAnd(input A, B, output Z);
  assign Z = A & B;
endmodule
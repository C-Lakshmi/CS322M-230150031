// XOR gate
module MyXor(input A, B, output Z);
  assign Z = A ^ B;
endmodule